
// zdf
module adder(
input wire a,
input wire b,
output wire c
);
asign c = a + b;
